`ifndef ADC_CONTROLLER_VH
`define ADC_CONTROLLER_VH
`define REG_ADC_CHANNEL_BYPASS_0 16'd0
`define REG_ADC_CHANNEL_BYPASS_1 16'd1
`define REG_ADC_CMON_EN          16'd2
`define REG_ADC_TMON_EN          16'd3
`define REG_ADC_EN               16'd4
`define REG_AVG_CONF             16'd5
`define REG_ADC_STATUS           16'd6
`endif
