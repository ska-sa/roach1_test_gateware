module TB_analogure_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
