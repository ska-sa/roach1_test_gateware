`ifndef POWER_MANAGER_VH
`define POWER_MANAGER_VH
`define REG_POWERSTATE        16'd0
`define REG_POWERUP           16'd1
`define REG_POWERDOWN         16'd2
`define REG_CRASH_CTRL        16'd3
`define REG_WATCHDOG_CTRL     16'd4
`define REG_WATCHDOG_CONF     16'd5
`define REG_CHS_SHUTDOWN_CTRL 16'd6
`define REG_ATXLOADRES_CTRL   16'd7
`define REG_PS_POWERGDS       16'd8
`endif
