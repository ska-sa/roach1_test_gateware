module qdr_controller(
  );
endmodule
