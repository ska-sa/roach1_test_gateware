module TB_sys_config();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
