module TB_iadc_controller();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
