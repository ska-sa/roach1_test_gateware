`timescale 1ns/10ps
`include "memlayout.v"
module gen_memlayout ();
  initial begin
    $display("#ifndef %s_%s_REGISTERS_H        ","`MODULE_ID","`REV_MAJOR");
    $display("#define %s_%s_REGISTERS_H        ","`MODULE_ID","`REV_MAJOR");
    $display("#define %s_FROM_BID_A        0x%x","`MODULE_ID",`FROM_BID_A);
    $display("#define %s_FROM_BID_L        0x%x","`MODULE_ID",`FROM_BID_L);
    $display("#define %s_FROM_REV_A        0x%x","`MODULE_ID",`FROM_REV_A);
    $display("#define %s_FROM_REV_L        0x%x","`MODULE_ID",`FROM_REV_L);
    $display("#define %s_FROM_LEVELS_A     0x%x","`MODULE_ID",`FROM_LEVELS_A);
    $display("#define %s_FROM_LEVELS_L     0x%x","`MODULE_ID",`FROM_LEVELS_L);
    $display("#define %s_FROM_ACMDATA_A    0x%x","`MODULE_ID",`FROM_ACMDATA_A);
    $display("#define %s_FROM_ACMDATA_L    0x%x","`MODULE_ID",`FROM_ACMDATA_L);
    $display("#define %s_ACM_AQUADS_A      0x%x","`MODULE_ID",`ACM_AQUADS_A);
    $display("#define %s_ACM_AQUADS_L      0x%x","`MODULE_ID",`ACM_AQUADS_L);
    $display("#define %s_ALC_FAULTVAL_A    0x%x","`MODULE_ID",`ALC_FAULTVAL_A);
    $display("#define %s_ALC_FAULTVAL_L    0x%x","`MODULE_ID",`ALC_FAULTVAL_L);
    $display("#define %s_ALC_HARDLEVEL_A   0x%x","`MODULE_ID",`ALC_HARDLEVEL_A);
    $display("#define %s_ALC_HARDLEVEL_L   0x%x","`MODULE_ID",`ALC_HARDLEVEL_L);
    $display("#define %s_ALC_SOFTLEVEL_A   0x%x","`MODULE_ID",`ALC_SOFTLEVEL_A);
    $display("#define %s_ALC_SOFTLEVEL_L   0x%x","`MODULE_ID",`ALC_SOFTLEVEL_L);
    $display("#define %s_ALC_ADCVAL_A      0x%x","`MODULE_ID",`ALC_ADC_VALUE_A);
    $display("#define %s_ALC_ADC_VALUE_L   0x%x","`MODULE_ID",`ALC_ADC_VALUE_L);
    $display("#define %s_ALC_RBUFF_A       0x%x","`MODULE_ID",`ALC_RBUFF_A);
    $display("#define %s_ALC_RBUFF_L       0x%x","`MODULE_ID",`ALC_RBUFF_L);
    $display("#define %s_PM_SHUTDOWN_A     0x%x","`MODULE_ID",`PC_SHUTDOWN_A);
    $display("#define %s_PM_SHUTDOWN_L     0x%x","`MODULE_ID",`PC_SHUTDOWN_L);
    $display("#define %s_PM_CHSALERT_A     0x%x","`MODULE_ID",`PC_CHASSIS_ALERT_A);
    $display("#define %s_PM_CHSALERT_L     0x%x","`MODULE_ID",`PC_CHASSIS_ALERT_L);
    $display("#define %s_PM_CRASH_A        0x%x","`MODULE_ID",`PC_CRASH_A);
    $display("#define %s_PM_CRASH_L        0x%x","`MODULE_ID",`PC_CRASH_L);
    $display("#define %s_PM_WATCHDOG_A     0x%x","`MODULE_ID",`PC_WATCHDOG_A);
    $display("#define %s_PM_WATCHDOG_L     0x%x","`MODULE_ID",`PC_WATCHDOG_L);
    $display("#define %s_PM_GA_A           0x%x","`MODULE_ID",`PC_GA_A);
    $display("#define %s_PM_GA_L           0x%x","`MODULE_ID",`PC_GA_L);
    $display("#define %s_PM_PD_A           0x%x","`MODULE_ID",`PC_PD_A);
    $display("#define %s_PM_PD_L           0x%x","`MODULE_ID",`PC_PD_L);
    $display("#define %s_PM_POWERUP_A      0x%x","`MODULE_ID",`PC_POWERUP_A);
    $display("#define %s_PM_POWERUP_L      0x%x","`MODULE_ID",`PC_POWERUP_L);
    $display("#define %s_IRQC_FLAG_A       0x%x","`MODULE_ID",`IRQC_FLAG_A);
    $display("#define %s_IRQC_FLAG_L       0x%x","`MODULE_ID",`IRQC_FLAG_L);
    $display("#define %s_IRQC_USER_A       0x%x","`MODULE_ID",`IRQC_USER_A);
    $display("#define %s_IRQC_USER_L       0x%x","`MODULE_ID",`IRQC_USER_L);
    $display("#define %s_IRQC_MASK_A       0x%x","`MODULE_ID",`IRQC_MASK_A);
    $display("#define %s_IRQC_MASK_L       0x%x","`MODULE_ID",`IRQC_MASK_L);
    $display("#define %s_BUSMON_ADDR_A     0x%x","`MODULE_ID",`BUSMON_ADDR_A);
    $display("#define %s_BUSMON_ADDR_L     0x%x","`MODULE_ID",`BUSMON_ADDR_L);
    $display("#define %s_BUSMON_CMND_A     0x%x","`MODULE_ID",`BUSMON_CMND_A);
    $display("#define %s_BUSMON_CMND_L     0x%x","`MODULE_ID",`BUSMON_CMND_L);
    $display("#define %s_BUSMON_DATA_A     0x%x","`MODULE_ID",`BUSMON_DATA_A);
    $display("#define %s_BUSMON_DATA_L     0x%x","`MODULE_ID",`BUSMON_DATA_L);
    $display("#define %s_BUSMON_COUNT_A    0x%x","`MODULE_ID",`BUSMON_COUNT_A);
    $display("#define %s_BUSMON_COUNT_L    0x%x","`MODULE_ID",`BUSMON_COUNT_L);
    $display("#define %s_BUSMON_CADDR_A    0x%x","`MODULE_ID",`BUSMON_CADDR_A);
    $display("#define %s_BUSMON_CADDR_L    0x%x","`MODULE_ID",`BUSMON_CADDR_L);
    $display("#define %s_BUSMON_CCMND_A    0x%x","`MODULE_ID",`BUSMON_CCMND_A);
    $display("#define %s_BUSMON_CCMND_L    0x%x","`MODULE_ID",`BUSMON_CCMND_L);
    $display("#define %s_BUSMON_CDATA_A    0x%x","`MODULE_ID",`BUSMON_CDATA_A);
    $display("#define %s_BUSMON_CDATA_L    0x%x","`MODULE_ID",`BUSMON_CDATA_L);
    $display("#define %s_BUSMON_OPCNT_A    0x%x","`MODULE_ID",`BUSMON_OPCNT_A);
    $display("#define %s_BUSMON_OPCNT_L    0x%x","`MODULE_ID",`BUSMON_OPCNT_L);
    $display("#define %s_AP_ADDR_A         0x%x","`MODULE_ID",`AP_ADDR_A);
    $display("#define %s_AP_ADDR_L         0x%x","`MODULE_ID",`AP_ADDR_L);
    $display("#define %s_AP_CMND_A         0x%x","`MODULE_ID",`AP_CMND_A);
    $display("#define %s_AP_CMND_L         0x%x","`MODULE_ID",`AP_CMND_L);
    $display("#define %s_FDBG_WCNT_A       0x%x","`MODULE_ID",`FLASH_DEBUG_WRITE_COUNT_A);
    $display("#define %s_FDBG_WCNT_L       0x%x","`MODULE_ID",`FLASH_DEBUG_WRITE_COUNT_L);
    $display("#define %s_FDBG_RCNT_A       0x%x","`MODULE_ID",`FLASH_DEBUG_READ_COUNT_A);
    $display("#define %s_FDBG_RCNT_L       0x%x","`MODULE_ID",`FLASH_DEBUG_READ_COUNT_L);
    $display("#define %s_FDBG_PCNT_A       0x%x","`MODULE_ID",`FLASH_DEBUG_PROG_COUNT_A);
    $display("#define %s_FDBG_PCNT_L       0x%x","`MODULE_ID",`FLASH_DEBUG_PROG_COUNT_L);
    $display("#define %s_FDBG_WFAILCNT_A   0x%x","`MODULE_ID",`FLASH_DEBUG_WRITE_FAIL_COUNT_A);
    $display("#define %s_FDBG_WFAILCNT_L   0x%x","`MODULE_ID",`FLASH_DEBUG_WRITE_FAIL_COUNT_L);
    $display("#define %s_FDBG_RFAILCNT_A   0x%x","`MODULE_ID",`FLASH_DEBUG_READ_FAIL_COUNT_A);
    $display("#define %s_FDBG_RFAILCNT_L   0x%x","`MODULE_ID",`FLASH_DEBUG_READ_FAIL_COUNT_L);
    $display("#define %s_FDBG_PFAILCNT_A   0x%x","`MODULE_ID",`FLASH_DEBUG_PROG_FAIL_COUNT_A);
    $display("#define %s_FDBG_PFAILCNT_L   0x%x","`MODULE_ID",`FLASH_DEBUG_PROG_FAIL_COUNT_L);
    $display("#define %s_FDBG_WTRANSCNT_A  0x%x","`MODULE_ID",`FLASH_DEBUG_WRITE_TRANS_COUNT_A);
    $display("#define %s_FDBG_WTRANSCNT_L  0x%x","`MODULE_ID",`FLASH_DEBUG_WRITE_TRANS_COUNT_L);
    $display("#define %s_FDBG_RTRANSCNT_A  0x%x","`MODULE_ID",`FLASH_DEBUG_READ_TRANS_COUNT_A);
    $display("#define %s_FDBG_RTRANSCNT_L  0x%x","`MODULE_ID",`FLASH_DEBUG_READ_TRANS_COUNT_L);
    $display("#define %s_FLASH_PAGESTAT_A  0x%x","`MODULE_ID",`FLASH_PAGE_STATUS_A);
    $display("#define %s_FLASH_PAGESTAT_L  0x%x","`MODULE_ID",`FLASH_PAGE_STATUS_L);
    $display("#define %s_FLASH_STATUS_A    0x%x","`MODULE_ID",`FLASH_STATUS_A);
    $display("#define %s_FLASH_STATUS_L    0x%x","`MODULE_ID",`FLASH_STATUS_L);
    $display("#define %s_FLASH_DPAGE_A     0x%x","`MODULE_ID",`FLASH_DIRTY_PAGE_A);
    $display("#define %s_FLASH_DPAGE_L     0x%x","`MODULE_ID",`FLASH_DIRTY_PAGE_L);
    $display("#define %s_FLASH_DATA_A      0x%x","`MODULE_ID",`FLASH_DATA_A);
    $display("#define %s_FLASH_DATA_L      0x%x","`MODULE_ID",`FLASH_DATA_L);
    $display("#endif");
    $finish;
  end
endmodule
