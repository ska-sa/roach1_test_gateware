`ifndef SYS_BLOCK_VH
`define SYS_BLOCK_VH
`define REG_BOARD_ID   3'd0
`define REG_REV_MAJOR  3'd1
`define REG_REV_MINOR  3'd2
`define REG_REV_RCS    3'd3
`define REG_SCRATCHPAD 3'd4
`endif
