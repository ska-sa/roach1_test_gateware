`ifndef BUS_MONITOR_VH
`define BUS_MONITOR_VH
`define REG_BUS_STATUS_0  16'd0
`define REG_BUS_STATUS_1  16'd1
`define REG_TIMEOUT_COUNT 16'd2
`define REG_MEMV_COUNT    16'd3
`define REG_UART_STATUS   16'd4
`endif
