`ifndef SYS_CONFIG_VH
`define SYS_CONFIG_VH
`define REG_BOARD_ID     16'd0
`define REG_REV_MAJOR    16'd1
`define REG_REV_MINOR    16'd2
`define REG_REV_RCS      16'd3
`define REG_RCS_UPTODATE 16'd4
`define REG_SYS_CONFIG   16'd5
`define REG_TIME_SEC_2   16'd6
`define REG_TIME_SEC_1   16'd7
`define REG_TIME_SEC_0   16'd8
`define REG_TIME_TICKER  16'd9
`endif
