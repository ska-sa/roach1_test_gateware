`ifndef DDR2_CPU_INTERFACE_VH
`define DDR2_CPU_INTERFACE_VH

`define REG_DDR2_PHY_READY 3'd0
`define REG_DDR2_SOFT_ADDR 3'd1
`define REG_DDR2_RESET     3'd2
`define REG_DDR2_BUS_RQST  3'd3
`define REG_DDR2_BUS_GRNTD 3'd4
`define REG_DDR2_FREQ      3'd5

`endif
