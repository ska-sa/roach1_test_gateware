module IBUF(
    I, O
  );
  input  I;
  output O;
endmodule
