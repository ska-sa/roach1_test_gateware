module iadc_test_harness(
  );
endmodule
