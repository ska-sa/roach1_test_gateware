module TB_v5c_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
