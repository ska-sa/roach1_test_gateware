module TB_misc();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
