module iadc_infrastructure(
  );
endmodule
