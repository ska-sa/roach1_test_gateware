module RAM4K9(
    RESET,
    CLKA,
    ADDRA11, ADDRA10, ADDRA9, ADDRA8, ADDRA7, ADDRA6, ADDRA5, ADDRA4, ADDRA3, ADDRA2, ADDRA1, ADDRA0,
    DINA8, DINA7, DINA6, DINA5,DINA4, DINA3, DINA2, DINA1, DINA0,
    DOUTA8, DOUTA7, DOUTA6, DOUTA5,DOUTA4, DOUTA3,DOUTA2,DOUTA1,DOUTA0,
    WIDTHA1, WIDTHA0, PIPEA, WMODEA, BLKA, WENA,
    CLKB,
    ADDRB11, ADDRB10, ADDRB9, ADDRB8, ADDRB7, ADDRB6, ADDRB5, ADDRB4, ADDRB3, ADDRB2, ADDRB1, ADDRB0,
    DINB8, DINB7, DINB6, DINB5,DINB4, DINB3, DINB2, DINB1, DINB0,
    DOUTB8, DOUTB7, DOUTB6, DOUTB5,DOUTB4, DOUTB3,DOUTB2,DOUTB1,DOUTB0,
    WIDTHB1, WIDTHB0, PIPEB, WMODEB, BLKB, WENB
  );
  input  RESET;
  input  CLKA;
  input  ADDRA11, ADDRA10, ADDRA9, ADDRA8, ADDRA7, ADDRA6, ADDRA5, ADDRA4, ADDRA3, ADDRA2, ADDRA1, ADDRA0;
  input  DINA8, DINA7, DINA6, DINA5,DINA4, DINA3, DINA2, DINA1, DINA0;
  output DOUTA8, DOUTA7, DOUTA6, DOUTA5,DOUTA4, DOUTA3,DOUTA2,DOUTA1,DOUTA0;
  input  WIDTHA1, WIDTHA0, PIPEA, WMODEA, BLKA, WENA;
  input  CLKB;
  input  ADDRB11, ADDRB10, ADDRB9, ADDRB8, ADDRB7, ADDRB6, ADDRB5, ADDRB4, ADDRB3, ADDRB2, ADDRB1, ADDRB0;
  input  DINB8, DINB7, DINB6, DINB5,DINB4, DINB3, DINB2, DINB1, DINB0;
  output DOUTB8, DOUTB7, DOUTB6, DOUTB5,DOUTB4, DOUTB3,DOUTB2,DOUTB1,DOUTB0;
  input  WIDTHB1, WIDTHB0, PIPEB, WMODEB, BLKB, WENB;
endmodule
