module TB_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
