module TB_qdr_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
