module TB_flashmem_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
