`ifndef RC_IRQ_CONTROLLER_H
`define RC_IRQ_CONTROLLER_H
`define REG_IRQC_FLAG 16'd0
`define REG_IRQC_USER 16'd1
`define REG_IRQC_MASK 16'd2
`endif
