module TB_xaui_fifo();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
