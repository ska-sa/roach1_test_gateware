`ifndef VALUE_STORAGE_VH
`define VALUE_STORAGE_VH
`define REG_RB_CTRL 16'd32
`endif
