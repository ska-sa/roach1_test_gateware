`ifndef DRAM_CPU_INTERFACE_VH
`define DRAM_CPU_INTERFACE_VH

`define REG_DRAM_PHY_READY 3'd0
`define REG_DRAM_RESET     3'd1
`define REG_DRAM_FREQ      3'd2

`endif
