module TB_ddr2_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
