module TB_epb_wb_bridge();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
