module TB_flashrom_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
