`ifndef CRC_VH
`define CRC_VH
`define CRC_ORDER 8
`define M_LENGTH  40

`define MESSAGE {1'b0,1'b1,6'd16,32'h0000_0000}
`define DIVISOR {7'b000_1001}
`endif
