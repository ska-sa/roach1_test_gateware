`ifndef SYS_BLOCK_VH
`define SYS_BLOCK_VH
`define REG_BOARD_ID     4'd0
`define REG_REV_MAJOR    4'd1
`define REG_REV_MINOR    4'd2
`define REG_REV_RCS      4'd3
`define REG_RCS_UPTODATE 4'd4
`define REG_SCRATCHPAD   4'd5
`define REG_SOFT_RESET   4'd6
`define REG_USER_IRQ     4'd7
`endif
