`ifndef VALUE_STORAGE_VH
`define VALUE_STORAGE_VH
`define REG_RB_CTRL      16'd32
`define REG_SAMPLE_COUNT 16'd33
`endif
