`ifndef DDR2_TEST_HARNESS_VH
`define DDR2_TEST_HARNESS_VH
`define REG_DDR2_TH_CTRL_0   5'd0
`define REG_DDR2_TH_CTRL_1   5'd1
`define REG_DDR2_TH_CTRL_2   5'd2
`define REG_DDR2_TH_CTRL_3   5'd3
`define REG_DDR2_TH_CTRL_4   5'd4
`endif
