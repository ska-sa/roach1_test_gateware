module TB_ddr2_cpu_interface();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
