module qdr_test_harness(
  );
endmodule
