`ifndef SYS_CONFIG_VH
`define SYS_CONFIG_VH
`define REG_BOARD_ID   16'd0
`define REG_REV_MAJOR  16'd1
`define REG_REV_MINOR  16'd2
`define REG_REV_RCS    16'd3
`define REG_SYS_CONFIG 16'd4
`endif
