module iadc_controller(
  );
endmodule
