module TB_qdr_cpu_interface();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
