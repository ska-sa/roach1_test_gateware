`timescale 1ns/1ps
module TB_fan_controller();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
