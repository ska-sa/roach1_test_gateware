module ddr2_cpu_interface(
  );
endmodule
