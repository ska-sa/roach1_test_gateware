module qdr_infrastructure(
  );
endmodule
