module BIBUF(
  D,E,Y,PAD
  );
  input D,E;
  output Y,PAD;
endmodule
