module qdr_cpu_interface(
  );
endmodule
