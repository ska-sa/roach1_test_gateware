module TB_lc_infrastructure();

  initial begin
    $display("PASSED");
    $finish;
  end

endmodule
