module ddr2_test_harness(
  );
endmodule
