`ifndef IADC_CONTROLLER_VH
`define IADC_CONTROLLER_VH

`define REG_IADC_RESET       4'd0 
`define REG_IADC_MODE        4'd1
`define REG_IADC_TWI_ADDR    4'd2
`define REG_IADC_TWI_DATA    4'd3
`define REG_IADC_TWI_TX      4'd4
`define REG_IADC_FIFODATA_4  4'd5
`define REG_IADC_FIFODATA_3  4'd6
`define REG_IADC_FIFODATA_2  4'd7
`define REG_IADC_FIFODATA_1  4'd8
`define REG_IADC_FIFODATA_0  4'd9
`define REG_IADC_FIFO_ADV    4'd10
`define REG_IADC_FIFO_STATUS 4'd11
`define REG_IADC_FIFO_CTRL   4'd12

`endif
