`ifndef QDR_CPU_INTERFACE_VH
`define QDR_CPU_INTERFACE_VH

`define REG_QDR_PHY_READY 3'd0
`define REG_QDR_RESET     3'd1

`endif
