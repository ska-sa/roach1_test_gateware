`ifndef DDR2_TEST_HARNESS_VH
`define DDR2_TEST_HARNESS_VH
`define REG_DDR2_TH_CTRL_0   7'd0
`define REG_DDR2_TH_CTRL_1   7'd1
`define REG_DDR2_TH_CTRL_2   7'd2
`define REG_DDR2_TH_CTRL_3   7'd3
`define REG_DDR2_TH_CTRL_4   7'd4
`define REG_DDR2_TH_CTRL_5   7'd5
`define REG_DDR2_TH_CTRL_6   7'd6
`endif
