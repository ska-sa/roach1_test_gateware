`ifndef XAUI_PIPE_VH 
`define XAUI_PIPE_VH

`define REG_TXDATA3        5'd0
`define REG_TXDATA2        5'd1
`define REG_TXDATA1        5'd2
`define REG_TXDATA0        5'd3
`define REG_TXADVANCE      5'd4
`define REG_TXSTATUS       5'd5
`define REG_RXDATA3        5'd6
`define REG_RXDATA2        5'd7
`define REG_RXDATA1        5'd8
`define REG_RXDATA0        5'd9
`define REG_RXADVANCE      5'd10
`define REG_RXSTATUS       5'd11
`define REG_LINKSTATUS     5'd12
`define REG_POWERDOWN      5'd13
`define REG_LOOPBACK       5'd14
`define REG_TXEN           5'd15
`define REG_RESET          5'd16
`define REG_RXPHYCONF      5'd17
`define REG_TXPHYCONF      5'd18
`define REG_UNUSED         5'd19

`endif
