module ddr2_infrastructure(
  );
endmodule
