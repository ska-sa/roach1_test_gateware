module qdrc_phy #(
    parameter DATA_WIDTH   = 18,
    parameter BW_WIDTH     = 2,
    parameter ADDR_WIDTH   = 21,
    parameter CLK_FREQ     = 200,
    parameter BURST_LENGTH = 4
  ) ( 
    input                       clk,
    input                       div_clk,
    input                       reset,
    output                      phy_rdy,
    output                      cal_fail,

    input                       phy_wr_strb,
    input    [ADDR_WIDTH - 1:0] phy_addr,

    input  [DATA_WIDTH*2 - 1:0] phy_wr_data,
    input    [BW_WIDTH*2 - 1:0] phy_wr_ben,

    input                       phy_rd_strb,
    output [DATA_WIDTH*2 - 1:0] phy_rd_data,

    output   [DATA_WIDTH - 1:0] qdr_d_rise,
    output   [DATA_WIDTH - 1:0] qdr_d_fall,
    input    [DATA_WIDTH - 1:0] qdr_q_rise,
    input    [DATA_WIDTH - 1:0] qdr_q_fall,

    output     [BW_WIDTH - 1:0] qdr_bw_n_rise,
    output     [BW_WIDTH - 1:0] qdr_bw_n_fall,
    output   [ADDR_WIDTH - 1:0] qdr_sa,
    output                      qdr_w_n,
    output                      qdr_r_n,

    output                      qdr_dll_off_n,

    output   [DATA_WIDTH - 1:0] dly_inc_dec_n,
    output   [DATA_WIDTH - 1:0] dly_en,
    output   [DATA_WIDTH - 1:0] dly_rst,

    input                       doffn,
    input                       cal_en,
    output                      cal_rdy,
    input                 [7:0] bit_select,
    input                       dll_en,
    input                       dll_inc_dec_n,
    input                       dll_rst,
    input                       align_strb,
    input                       align_en,
    output                [1:0] data_value,
    output                      data_sampled,
    output                      data_valid
  );

  reg cal_en_R;
  reg cal_en_RR;

  always @(posedge clk) begin
    cal_en_R  <= cal_en;
    cal_en_RR <= cal_en_R;
  end

  assign cal_fail = 1'b0;
  assign phy_rdy  = !cal_en_RR;

  wire cal_busy = cal_en_RR;
  wire cal_w_n;
  wire cal_r_n;
  wire [DATA_WIDTH - 1:0] cal_qdr_q_fall;
  wire [DATA_WIDTH - 1:0] cal_qdr_q_rise;

  assign qdr_d_rise = cal_busy ? {DATA_WIDTH{1'b1}} : phy_wr_data[DATA_WIDTH - 1:0];
  assign qdr_d_fall = cal_busy ? {DATA_WIDTH{1'b0}} : phy_wr_data[2*DATA_WIDTH - 1:DATA_WIDTH];

  assign qdr_bw_n_rise = cal_busy ? {BW_WIDTH{1'b0}} : ~phy_wr_ben[BW_WIDTH - 1:0];
  assign qdr_bw_n_fall = cal_busy ? {BW_WIDTH{1'b0}} : ~phy_wr_ben[BW_WIDTH*2 - 1:BW_WIDTH];

  assign qdr_sa = cal_busy ? {ADDR_WIDTH{1'b0}} : phy_addr;

  assign qdr_w_n = cal_busy ? cal_w_n : !phy_wr_strb;
  assign qdr_r_n = cal_busy ? cal_r_n : !phy_rd_strb;

  assign phy_rd_data = {cal_qdr_q_fall, cal_qdr_q_rise};

  /* cal sm */
  reg [1:0] state;
  localparam STATE_IDLE  = 2'd0;
  localparam STATE_WRITE = 2'd1;
  localparam STATE_READ  = 2'd2;

  always @(posedge clk) begin
    if (reset) begin
      state <= STATE_IDLE;
    end else begin
      case (state)
        STATE_IDLE: begin
          if (cal_busy) 
            state <= STATE_WRITE;
        end
        STATE_WRITE: begin
          state <= STATE_READ;
        end
        STATE_READ: begin
        end
      endcase
    end

    if (!cal_busy) 
      state <= STATE_IDLE;
  end

  assign cal_w_n = state == STATE_WRITE ? 1'b0 : 1'b1;
  assign cal_r_n = state == STATE_READ  ? 1'b0 : 1'b1;

  reg cal_rdyR;
  reg cal_rdyRR;
  always @(posedge div_clk) begin
    cal_rdyR  <= state == STATE_READ;
    cal_rdyRR <= cal_rdyR;
  end
  assign cal_rdy = cal_rdyRR;

  /* bit align */

  qdrc_phy_train #(
    .DATA_WIDTH (DATA_WIDTH)
  ) qdrc_phy_train_inst (
    .clk           (div_clk),
    .q_rise        (qdr_q_rise),
    .q_fall        (qdr_q_fall),
    .dly_inc_dec_n (dly_inc_dec_n),
    .dly_en        (dly_en),
    .dly_rst       (dly_rst),
    .bit_select    (bit_select),
    .dll_en        (dll_en),
    .dll_inc_dec_n (dll_inc_dec_n),
    .dll_rst       (dll_rst),
    .data_value    (data_value),
    .data_sampled  (data_sampled),
    .data_valid    (data_valid)    
  );

  qdrc_phy_align #(
    .DATA_WIDTH (DATA_WIDTH)
  ) qdrc_phy_align_inst (
    .clk           (clk),
    .divclk        (div_clk),
    .bit_select    (bit_select),
    .align_strb    (align_strb),
    .align_en      (align_en),
    .q_rise        (qdr_q_rise),
    .q_fall        (qdr_q_fall),
    .cal_rise      (cal_qdr_q_rise),
    .cal_fall      (cal_qdr_q_fall)
  );
  assign qdr_dll_off_n = doffn;
endmodule
