module TB_xaui_pipe();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
