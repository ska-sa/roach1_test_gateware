module TB_ten_gig_eth();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
