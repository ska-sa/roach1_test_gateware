module TB_qdr_controller();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
