module TB_iadc_infrastructure();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
