module TB_toplevel();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule
