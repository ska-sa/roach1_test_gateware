`ifndef DDR2_TEST_HARNESS_VH
`define DDR2_TEST_HARNESS_VH
`define REG_DDR2_TH_CTRL_0   4'd0
`define REG_DDR2_TH_CTRL_1   4'd1
`define REG_DDR2_TH_CTRL_2   4'd2
`endif
