`ifndef LEVEL_CHECKER_VH
`define LEVEL_CHECKER_VH
`define REG_SOFT_THRESH_VALID 16'h80
`define REG_HARD_THRESH_VALID 16'h81
`define REG_SOFT_VIOL_SOURCE  16'h82
`define REG_SOFT_VIOL_VALUE   16'h83
`define REG_HARD_VIOL_SOURCE  16'h84
`define REG_HARD_VIOL_VALUE   16'h85
`define REG_VINRANGE_0        16'h86
`define REG_VINRANGE_1        16'h87
`endif
