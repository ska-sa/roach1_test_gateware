`ifndef XAUI_PIPE_MEM_H 
`define XAUI_PIPE_MEM_H

`define XAUI_TXDATA_A         6'd0
`define XAUI_TXSTATUS_A       6'd1
`define XAUI_RXDATA_A         6'd2
`define XAUI_RXSTATUS_A       6'd3
`define XAUI_LINKSTATUS_A     6'd4
`define XAUI_LOOPBACK_A       6'd5
`define XAUI_TXEN_A           6'd6
`define XAUI_RESET_A          6'd7
`define XAUI_SRESET_A         6'd8
`define XAUI_POWERDOWN_A      6'd9

`define XAUI_MGT_STATUS_0_A   6'd10
`define XAUI_MGT_STATUS_1_A   6'd11
`define XAUI_MGT_PDIFF_A      6'd12
`define XAUI_MGT_CBSKEW_A     6'd13

`define XAUI_MGT_CHBOND_ERRORS_0_A      6'd14
`define XAUI_MGT_CHBOND_ERRORS_1_A      6'd15
`define XAUI_MGT_CHBOND_ERRORS_2_A      6'd16
`define XAUI_MGT_CHBOND_ERRORS_3_A      6'd17

`define XAUI_MGT_CLK_CORR_ERRORS_0_A    6'd18
`define XAUI_MGT_CLK_CORR_ERRORS_1_A    6'd19
`define XAUI_MGT_CLK_CORR_ERRORS_2_A    6'd20
`define XAUI_MGT_CLK_CORR_ERRORS_3_A    6'd21

`define XAUI_MGT_CLK_CORR_EVENTS_0_A    6'd22
`define XAUI_MGT_CLK_CORR_EVENTS_1_A    6'd23
`define XAUI_MGT_CLK_CORR_EVENTS_2_A    6'd24
`define XAUI_MGT_CLK_CORR_EVENTS_3_A    6'd25

`define XAUI_MGT_CHBOND_EVENTS_0_A    6'd26
`define XAUI_MGT_CHBOND_EVENTS_1_A    6'd27
`define XAUI_MGT_CHBOND_EVENTS_2_A    6'd28
`define XAUI_MGT_CHBOND_EVENTS_3_A    6'd29

`endif
