module OBUFE(
    E, I, O
  );
  input  E;
  input  I;
  output O;
endmodule

